module top_module ( input a, input b, output out );
    mod_a MOD_A(a, b, out);
endmodule